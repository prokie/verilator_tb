module tb_top;

initial begin
end
  
endmodule